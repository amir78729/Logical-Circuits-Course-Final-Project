`timescale 1ns / 1ps
`default_nettype none

/*
**********************************************************
** Logic Design Final Project Fall, 2'b10019 Semester
** Amirkabir University of Technology (Tehran Polytechnic)
** Department of Computer Engineering (CEIT-AUT)
** Logic Circuit Design Laboratory
** https://ceit.aut.ac.ir
**********************************************************
** Student ID: 9731078 (Negin HajiSobhani)
** Student ID: 9731096 (Amirhossein Alibakhshi)
**********************************************************
** Module Name: LogicHealthcareSystemController
**********************************************************
** Additional Comments:
*/

module LogicHealthcareSystemController(  
    clock,
    presureAbnormality,
    bloodAbnormality,
    fallDetected,
    temperatureAbnormality,
    nervousAbnormality,
    abnormaliryWarning);
  
input clock;
input presureAbnormality;
input bloodAbnormality;
input fallDetected;
input temperatureAbnormality;
input [1:0] nervousAbnormality;
output reg [2:0] abnormaliryWarning;

	///////////// FULLADDER VERSION /////////////
	/*
	Additional comments:
	
	At first we concatinate our 6 inputs into a 6digit
	binary string(serial!)
	
	serial:
	 _____________________________________
    |     |     |     |     |     |     |
    |  5  |  4  |  3  |  2  |  1  |  0  |
    |_____|_____|_____|_____|_____|_____|
	 
	 Then we seperate "serial" into 3 equal parts:
	 _____________ _____________ _____________
    |     |     | |     |     | |     |     |
    |  5  |  4  | |  3  |  2  | |  1  |  0  |
    |_____|_____| |_____|_____| |_____|_____|
	 
	 
			_____________ 
			|     |     |  
    each	|  X  |  Y  | has 3 different moods:
			|_____|_____|
	
	1) "0" (00) one,
	2) "1" (01) one, and
	3) "2" (10) one
	
	the 2bit number in paranthesize is number of ones in each
	part that can be generated by:  " { X and Y , X xor Y } "
	because of this table:
	
	X   Y     A(XandY)   B(XxorY)    decimal
	0   0         0          0        0 (00)
	0   1         0          1        1 (01)
	1   0         0          1        1 (01)
	1   1         1          0        2 (11)
	
	by adding this numbers together (by using fullAdders) we can
	calculate number of ones in "serial" :)
	*/
	wire [5:0] serial;
	assign serial = {presureAbnormality, bloodAbnormality, fallDetected, temperatureAbnormality, nervousAbnormality[0], nervousAbnormality[1]};
	wire [2:0] result;
	wire [2:0] a, b, r;
	wire middleCarry1, temp1, temp2, temp3;
	
	and a2(a[2], serial[5], serial[4]);
	xor b2(b[2], serial[5], serial[4]);
	
	and a1(a[1], serial[3], serial[2]);
	xor b1(b[1], serial[3], serial[2]);
	
	and a0(a[0], serial[1], serial[0]);
	xor b0(b[0], serial[1], serial[0]);
	
	fullAdder f0(b[2], b[1], 1'b0, r[0], middleCarry1);
	fullAdder f1(a[2], a[1], middleCarry1, r[1], r[2]);
	
	fullAdder F0(b[0], r[0], 1'b0, result[0], temp1);
	fullAdder F1(a[0], r[1], temp1, result[1], temp2);
	fullAdder F2(1'b0, r[2], temp2, result[2], temp3);
	
	//output :
	always @ (posedge clock)begin
		assign abnormaliryWarning = result;
	end





	/*
	///////////// MOORE MACHINE CONCAT VERSION /////////////
	//Additional comments:
	//If the inputs change during the programming, the serial is not
	//going to change!
	
   //concatinating inputs :
	wire [5:0] serial;
	assign serial = {presureAbnormality, bloodAbnormality, fallDetected, temperatureAbnormality, nervousAbnormality[0], nervousAbnormality[1]};
	//states definition :
	parameter
		S0 = 3'b000,// no "1" enserted
		S1 = 3'b001,// 1 "1" enserted
		S2 = 3'b010,// 2 "1"s enserted
		S3 = 3'b011,// 3 "1"s enserted
		S4 = 3'b100,// 4 "1"s enserted
		S5 = 3'b101,// 5 "1"s enserted
		S6 = 3'b110;// 6 "1"s enserted
	reg [2:0] state = S0;	
	integer i = 0;
	// the bit we are controling in each clock
	wire x = serial[i];
	//next states:
	always @ (posedge clock ) begin
		case(state)
			S0:
			begin 
				if (x) begin 
					state = S1;
					$monitor ("-------------------------\n%d error founded!", state);
				end
				i = i + 1;
			end
			S1:
			begin 
				if (x) begin 
					state = S2;
					$monitor ("-------------------------\n%d errors founded!", state);
				end
				i = i + 1;
			end
			S2:
			begin 
				if (x) begin 
					state = S3;
					$monitor ("-------------------------\n%d errors founded!", state);
				end
				i = i + 1;
			end
			S3:
			begin 
				if (x) begin 
					state = S4;
					$monitor ("-------------------------\n%d errors founded!", state);
				end
				i = i + 1;
			end
			S4:
			begin 
				if (x) begin 
					state = S5;
					$monitor ("-------------------------\n%d errors founded!", state);
				end
				i = i + 1;
			end
			S5:
			begin 
				if (x) begin 
					state = S6;
					$monitor ("-------------------------\n%d errors founded!", state);
				end
			end
			S6: ;
		endcase
		//assign abnormaliryWarning = presureAbnormality+ bloodAbnormality+ fallDetected+ temperatureAbnormality+ nervousAbnormality[0]+ nervousAbnormality[1];
	end
	always @ (posedge clock)begin
		assign abnormaliryWarning = state;
	end
	*/
	
	
	
	
	
	/*
	///////////// SUM VERSION /////////////
	//Additional comments:
	//for testing in testbenchs
	
	
	wire [2:0] sum = presureAbnormality+ bloodAbnormality+ fallDetected+ temperatureAbnormality+ nervousAbnormality[0]+ nervousAbnormality[1];
	//output :
	always @ (posedge clock)begin
		assign abnormaliryWarning = sum;
	end
	*/
	
	
	
endmodule
